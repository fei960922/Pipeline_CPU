/*
	
	  Computer System (1) ------ Final Project
		MIPS 5-Level Pipeline CPU (Advanced)

		Author: 	Xu Yifei	&	Zhang Yiyi
		Stu. ID:	5130309056	&	5132409031
		Class: 		F1324004(ACM2013)
		College:	Zhiyuan College
		University: Shanghai Jiao Tong University

		File type:	Verilog --- Test
		File name:	Final Test
		
*/

`include "pipeline.v"

module final_test;

endmodule